`define no_of_frames 1
